module dom_conv #()(  
  input                                      valid_o,
  input                                      wt_o,
  input                  [I_FDSSI_WIDTH-1:0] FDSSI_o,
  input                  [FIFO_NUM_O_BLK-1:0] FDSTI_o_all,
  input                    [I_SSI_WIDTH-1:0] SSI_o,
  input                   [I_SAM_OFFSET-1:0] s_o,
  input                                       ready_o,
  input                   [I_DATA_WIDTH-1:0]  data_o
  );


endmodule